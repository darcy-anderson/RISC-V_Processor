`timescale 1ns / 1ps

module instr_mem(
	input clk,
  input [31:0] pc_addr, // Input address from program counter
  output [31:0] instr_out
);

  (* ram_style = "block" *) reg [31:0] instr_rom [511:0];
  reg [31:0] instr_read;

  initial $readmemh("main.mem", instr_rom);

	always @(posedge clk) instr_read = instr_rom[pc_addr[12:2]];

  assign instr_out = instr_read;

endmodule